-- tb_RCA.vhd : testbench
library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
entity tb_RCA is
end entity tb_RCA;
